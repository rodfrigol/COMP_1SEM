library verilog;
use verilog.vl_types.all;
entity q53 is
    port(
        Si              : out    vl_logic;
        Ai              : in     vl_logic;
        Eimenos1        : in     vl_logic;
        Bi              : in     vl_logic;
        Ei              : out    vl_logic
    );
end q53;
