library verilog;
use verilog.vl_types.all;
entity b3 is
    port(
        F               : out    vl_logic;
        c               : in     vl_logic;
        d               : in     vl_logic;
        a               : in     vl_logic;
        b               : in     vl_logic
    );
end b3;
