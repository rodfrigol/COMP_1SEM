library verilog;
use verilog.vl_types.all;
entity q5_vlg_vec_tst is
end q5_vlg_vec_tst;
