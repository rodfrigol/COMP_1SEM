library verilog;
use verilog.vl_types.all;
entity b3_vlg_vec_tst is
end b3_vlg_vec_tst;
