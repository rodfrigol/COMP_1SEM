library verilog;
use verilog.vl_types.all;
entity q43_vlg_check_tst is
    port(
        F               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end q43_vlg_check_tst;
