library verilog;
use verilog.vl_types.all;
entity q53final is
    port(
        F8              : out    vl_logic;
        M               : in     vl_logic;
        S1              : in     vl_logic;
        S0              : in     vl_logic;
        Cin             : in     vl_logic;
        A1              : in     vl_logic;
        B1              : in     vl_logic;
        A2              : in     vl_logic;
        B2              : in     vl_logic;
        A3              : in     vl_logic;
        B3              : in     vl_logic;
        A4              : in     vl_logic;
        B4              : in     vl_logic;
        A5              : in     vl_logic;
        B5              : in     vl_logic;
        A6              : in     vl_logic;
        B6              : in     vl_logic;
        A7              : in     vl_logic;
        B7              : in     vl_logic;
        A8              : in     vl_logic;
        B8              : in     vl_logic;
        F1              : out    vl_logic;
        F2              : out    vl_logic;
        F3              : out    vl_logic;
        F4              : out    vl_logic;
        F5              : out    vl_logic;
        F6              : out    vl_logic;
        F7              : out    vl_logic;
        Cout            : out    vl_logic
    );
end q53final;
