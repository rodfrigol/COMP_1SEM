library verilog;
use verilog.vl_types.all;
entity b3_vlg_check_tst is
    port(
        F               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end b3_vlg_check_tst;
