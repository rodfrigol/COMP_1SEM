library verilog;
use verilog.vl_types.all;
entity q53_vlg_check_tst is
    port(
        Ei              : in     vl_logic;
        Si              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end q53_vlg_check_tst;
