library verilog;
use verilog.vl_types.all;
entity q53_vlg_check_tst is
    port(
        Fi              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end q53_vlg_check_tst;
