library verilog;
use verilog.vl_types.all;
entity q62_vlg_check_tst is
    port(
        C0              : in     vl_logic;
        M1              : in     vl_logic;
        M2              : in     vl_logic;
        M3              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end q62_vlg_check_tst;
