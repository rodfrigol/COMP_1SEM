library verilog;
use verilog.vl_types.all;
entity q52_vlg_check_tst is
    port(
        Y1imenos1       : in     vl_logic;
        Y3imenos1       : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end q52_vlg_check_tst;
