library verilog;
use verilog.vl_types.all;
entity q52_vlg_check_tst is
    port(
        Q1              : in     vl_logic;
        Q2              : in     vl_logic;
        Q3              : in     vl_logic;
        Q4              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end q52_vlg_check_tst;
