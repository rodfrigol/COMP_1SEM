library verilog;
use verilog.vl_types.all;
entity q53final_vlg_vec_tst is
end q53final_vlg_vec_tst;
