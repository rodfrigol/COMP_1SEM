library verilog;
use verilog.vl_types.all;
entity q62 is
    port(
        C0              : out    vl_logic;
        A0              : in     vl_logic;
        B0              : in     vl_logic;
        M1              : out    vl_logic;
        A1              : in     vl_logic;
        B1              : in     vl_logic;
        M2              : out    vl_logic;
        M3              : out    vl_logic
    );
end q62;
