library verilog;
use verilog.vl_types.all;
entity q61_vlg_check_tst is
    port(
        C               : in     vl_logic;
        F               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end q61_vlg_check_tst;
