library verilog;
use verilog.vl_types.all;
entity q51_vlg_sample_tst is
    port(
        X0              : in     vl_logic;
        X1              : in     vl_logic;
        X2              : in     vl_logic;
        X3              : in     vl_logic;
        X4              : in     vl_logic;
        X5              : in     vl_logic;
        X6              : in     vl_logic;
        X7              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end q51_vlg_sample_tst;
