library verilog;
use verilog.vl_types.all;
entity q4_vlg_vec_tst is
end q4_vlg_vec_tst;
