library verilog;
use verilog.vl_types.all;
entity q53_vlg_vec_tst is
end q53_vlg_vec_tst;
