library verilog;
use verilog.vl_types.all;
entity q43_vlg_vec_tst is
end q43_vlg_vec_tst;
