library verilog;
use verilog.vl_types.all;
entity q61 is
    port(
        F               : out    vl_logic;
        S1              : in     vl_logic;
        A               : in     vl_logic;
        C0              : in     vl_logic;
        B               : in     vl_logic;
        M               : in     vl_logic;
        S0              : in     vl_logic;
        C               : out    vl_logic
    );
end q61;
