library verilog;
use verilog.vl_types.all;
entity q52_vlg_vec_tst is
end q52_vlg_vec_tst;
