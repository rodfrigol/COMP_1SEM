library verilog;
use verilog.vl_types.all;
entity q42_vlg_check_tst is
    port(
        Z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end q42_vlg_check_tst;
