library verilog;
use verilog.vl_types.all;
entity q52 is
    port(
        Y1imenos1       : out    vl_logic;
        Y1i             : in     vl_logic;
        Y3i             : in     vl_logic;
        Ai              : in     vl_logic;
        Bi              : in     vl_logic;
        Y3imenos1       : out    vl_logic
    );
end q52;
