library verilog;
use verilog.vl_types.all;
entity lab1 is
    port(
        f               : out    vl_logic;
        X3              : in     vl_logic;
        X2              : in     vl_logic;
        X1              : in     vl_logic;
        X0              : in     vl_logic
    );
end lab1;
