library verilog;
use verilog.vl_types.all;
entity q53final_vlg_check_tst is
    port(
        Cout            : in     vl_logic;
        F1              : in     vl_logic;
        F2              : in     vl_logic;
        F3              : in     vl_logic;
        F4              : in     vl_logic;
        F5              : in     vl_logic;
        F6              : in     vl_logic;
        F7              : in     vl_logic;
        F8              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end q53final_vlg_check_tst;
