library verilog;
use verilog.vl_types.all;
entity q5_vlg_check_tst is
    port(
        A               : in     vl_logic;
        Y0              : in     vl_logic;
        Y1              : in     vl_logic;
        Y2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end q5_vlg_check_tst;
