library verilog;
use verilog.vl_types.all;
entity q51 is
    port(
        A               : out    vl_logic;
        X4              : in     vl_logic;
        X6              : in     vl_logic;
        X7              : in     vl_logic;
        X5              : in     vl_logic;
        X0              : in     vl_logic;
        X2              : in     vl_logic;
        X3              : in     vl_logic;
        X1              : in     vl_logic;
        Y2              : out    vl_logic;
        Y1              : out    vl_logic;
        Y0              : out    vl_logic
    );
end q51;
