library verilog;
use verilog.vl_types.all;
entity q62_vlg_vec_tst is
end q62_vlg_vec_tst;
