library verilog;
use verilog.vl_types.all;
entity q51_vlg_vec_tst is
end q51_vlg_vec_tst;
