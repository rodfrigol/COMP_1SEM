library verilog;
use verilog.vl_types.all;
entity q61_vlg_vec_tst is
end q61_vlg_vec_tst;
