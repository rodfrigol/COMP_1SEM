library verilog;
use verilog.vl_types.all;
entity q51 is
    port(
        F               : out    vl_logic;
        B               : in     vl_logic;
        A               : in     vl_logic
    );
end q51;
