library verilog;
use verilog.vl_types.all;
entity q42_vlg_vec_tst is
end q42_vlg_vec_tst;
