library verilog;
use verilog.vl_types.all;
entity questao611_vlg_vec_tst is
end questao611_vlg_vec_tst;
