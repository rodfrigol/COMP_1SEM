library verilog;
use verilog.vl_types.all;
entity Block2 is
    port(
        y               : out    vl_logic;
        S0              : in     vl_logic;
        X0              : in     vl_logic;
        X1              : in     vl_logic;
        S1              : in     vl_logic;
        X2              : in     vl_logic;
        X3              : in     vl_logic
    );
end Block2;
