library verilog;
use verilog.vl_types.all;
entity q53 is
    port(
        Fi              : out    vl_logic;
        M               : in     vl_logic;
        Ai              : in     vl_logic;
        S0              : in     vl_logic;
        Bi              : in     vl_logic;
        S1              : in     vl_logic;
        Cin             : in     vl_logic
    );
end q53;
